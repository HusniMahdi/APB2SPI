package apb_agent_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::* ;
	import test_param_pkg::* ;
	
	`include "apb_seq_item.sv"
	`include "apb_driver_proxy.sv"
	`include "apb_monitor.sv"
	`include "apb_sqncr.sv"
	`include "apb_cov.sv"
	`include "apb_agent_config.sv"
	`include "apb_agent.sv"

        
endpackage 
